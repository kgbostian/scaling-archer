----------------------------------------------------------------------------------
-- Mojo_top VHDL
-- Translated from Mojo-base Verilog project @ http://embeddedmicro.com/frontend/files/userfiles/files/Mojo-Base.zip
-- by Xark
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity mojo_top is
	port (
		clk					: in  std_logic;		-- 50Mhz clock
		rst_n					: in  std_logic;		-- "reset" button input (negative logic)
		cclk					: in  std_logic;		-- configuration clock (?) from AVR (to detect when AVR ready)
		--led					: out std_logic_vector(7 downto 0);	 -- 8 LEDs on Mojo board
		--Anode Mux
		data_in  			: in std_logic_vector(3 downto 0);
		data_out_mux 		: out std_logic_vector(15 downto 0);
		--Decoder
		data_out_decoder	: out std_logic_vector(3 downto 0);
		--Counter "Clock" signal
		counter_clock		: in std_logic -- generated by RPI
		
	);
end mojo_top;

architecture RTL of mojo_top is

signal rst	       : std_logic;     -- reset signal (rst_n inverted for postive logic)
--Mux selector pins (bit 0,1), Decoder selector pins (bit 2,3)
signal sel             : std_logic_vector(3 downto 0);
signal out_mux_latch   : std_logic_vector(15 downto 0);
--RPI code needs to be modified to set write to the next line that is to be displayed


begin
--rst <= not rst_n;
--led <= "10000000" when sel = "00" else
--		 "01000000" when sel = "01" else
--		 "00100000" when sel = "10" else
--		 "00010000" when sel = "11" else
--		 "00000000";


-- Bus multiplexer (anode side)
--data_out_mux <= data_in & "000000000000" when sel(1 downto 0) = "00" else
--				  "0000" & data_in & "00000000" when sel(1 downto 0) = "01" else
--                "00000000" & data_in & "0000" when sel(1 downto 0) = "10" else
--				  "000000000000" & data_in when sel(1 downto 0) = "11" else
--               (others => '0');

--Counter
process (counter_clock, rst_n) --Counter clock and reset button sensitivity list
begin

--reset
if(rst_n = '0') then 
	sel <= "0000";
	data_out_mux <= (others => '0');
	out_mux_count <= 0;
--counter inc
elsif(counter_clock'event and counter_clock = '1') then
	sel <= sel + 1;
	out_latch_count <= out_latch_count+1;
	if(sel(1 downto 0) = "00") then
	    out_mux_latch(3 downto 0) <= data_in;
	elsif(sel(1 downto 0) = "01") then
	    out_mux_latch(7 downto 4) <= data_in;
	elsif(sel(1 downto 0) = "10") then
	    out_mux_latch(11 downto 8) <= data_in;
	elsif(sel(1 downto 0) = "11") then
	    out_mux_latch(15 downto 12 <= data_in;
	    data_out_mux <= out_mux_latch;
	else
	    data_out_mux <= (others => '0');
	end if;
end if;
end process;


--Decoder
--sel(3 downto 2)
data_out_decoder <= "1000" when sel(3 downto 2) = "00" else
                    "0001" when sel(3 downto 2) = "01" else
                    "0010" when sel(3 downto 2) = "10" else
                    "0100" when sel(3 downto 2) = "11" else
                    (others => '0');

end RTL;
